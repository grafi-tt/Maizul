library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.types.all;

-- currently, BlockRAM is merely ROM

entity BlkRAM is
    port (
        clk : in std_logic;
        addr : in blkram_addr;
        instruction : out instruction_t := (others => '0'));
end entity;

architecture instance of BlkRAM is
    type blkram_t is array (0 to 31) of instruction_t;
    signal RAM : blkram_t := (
        "00010100000000010000000000100000", -- r1 = r0 | 32
        "10000100010000100000000000000000", -- mem(r2) = r2
        "00000000010000100000000000000001", -- r2 = r2 + 1
        "00000100001000010000000000000001", -- r1 = r1 - 1
        "11000100001000000000000000000001", -- jmp to inst1 if r1 != 0
        "01001000010000000000000000000001", -- print r2, which should be 32
        "00000100010000100000000000000100", -- r2 = r2 - 4
        "10000000010000110000000000000000", -- r3 = mem(r2)
        "10000000010001000000000000000001", -- r4 = mem(r2+1word)
        "10000000010001010000000000000010", -- r5 = mem(r2+2word)
        "10000000010001100000000000000011", -- r6 = mem(r2+3word)
        "01001000110000000000000000000001", -- print r6
        "01001000101000000000000000000001", -- print r5
        "01001000100000000000000000000001", -- print r4
        "01001000011000000000000000000001", -- print r3
        "11000100010000000000000000000110", -- jmp to inst6 if r2 != 0
        "01010000000000000000000000010000", -- jmp to myself (halt)
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000"
    );

begin
    everyClock : process(clk)
    begin
        if (rising_edge(clk)) then
            instruction <= RAM(to_integer(unsigned(addr(4 downto 0))));
        end if;
    end process;

end architecture;
