library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.types.all;

-- currently, BlockRAM is merely ROM

entity BlkRAM is
    port (
        clk : in std_logic;
        addr : in blkram_addr;
        instruction : out instruction_t := (others => '0'));
end entity;

architecture instance of BlkRAM is
    type blkram_t is array (0 to 31) of instruction_t;
    signal RAM : blkram_t := (
        "00010100000000100000000000101000", -- r2 = r0 | 40
        "01010100000111110000000000000100", -- r31 = nextPC, jmp to inst4:fib
        "01001000001000000000000000000001", -- print r1
        "01010000000000000000000000000011", -- halt
        "00001100010000110000000000000010", -- r3 = r2 < 2
        "00010100000000010000000000000001", -- r1 = r0 | 1
        "11000100011000000000000000010100", -- jmp to inst20:fibret if r3 != 0
        "00000011110111100000000000001000", -- r30 = r30 + 8
        "10000111110111111111111111111110", -- mem(r30 - 2word) = r31
        "10000111110000101111111111111111", -- mem(r30 - 1word) = r2
        "00000100010000100000000000000001", -- r2 = r2 - 1
        "01010100000111110000000000000100", -- r31 = nextPC, jmp to inst4:fib
        "10000011110000101111111111111111", -- r2 = mem(r30 - 1word)
        "10000111110000011111111111111111", -- mem(r30 - 1word) = r1
        "00000100010000100000000000000010", -- r2 = r2 - 2
        "01010100000111110000000000000100", -- r31 = nextPC, jmp to inst4:fib
        "10000011110000101111111111111111", -- r2 = mem(r30 - 1word)
        "01000000001000100000100000000000", -- r1 = r1 + r2
        "10000011110111111111111111111110", -- r31 = mem(r30 - 2word)
        "00000111110111100000000000001000", -- r30 = r30 - 8
        "01011011111000000000000000000000", -- r0 = nextPC, jmp to r31
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000"
    );

begin
    everyClock : process(clk)
    begin
        if (rising_edge(clk)) then
            instruction <= RAM(to_integer(unsigned(addr(4 downto 0))));
        end if;
    end process;

end instance;
