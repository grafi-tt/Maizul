library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.types.all;

-- currently, BlockRAM is merely ROM

entity BlkRAM is
    port (
        clk : in std_logic;
        addr : in blkram_addr;
        instruction : out instruction_t := (others => '0'));
end entity;

architecture instance of BlkRAM is
    type blkram_t is array (0 to 31) of instruction_t;
    signal RAM : blkram_t := (
        "00010100000111100000000000000000",
        "00101000000111010000000000001100",
        "00010100000000100000000000001010", -- fib 10
        "01010100000111110000000000000110",
        "01011100001000000000000000000001",
        "01010000000000000000000000000101",
        "00001100010000110000000000000010",
        "00010100000000010000000000000001",
        "10000100011000000000000000010110",
        "00000011101111010000000000000010",
        "01001111101111111111111111111110",
        "01001111101000101111111111111111",
        "00000100010000100000000000000001",
        "01010100000111110000000000000110",
        "01001011101000101111111111111111",
        "01001111101000011111111111111111",
        "00000100010000100000000000000010",
        "01010100000111110000000000000110",
        "01001011101000101111111111111111",
        "01000000001000100000100000000000",
        "01001011101111111111111111111110",
        "00000111101111010000000000000010",
        "01011011111000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000"
    );

begin
    everyClock : process(clk)
    begin
        if (rising_edge(clk)) then
            instruction <= RAM(to_integer(unsigned(addr(4 downto 0))));
        end if;
    end process;

end instance;
